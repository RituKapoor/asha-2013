  8 u � � � &Laddar ned aktiverare: %0U kB / %1U kB ;Något blev fel vid uppdateringen av meddelande­aktivering (Du måste uppdatera meddelandeaktivering !Uppdaterar meddelande­aktivering 6Minnet fullt. Radera några filer för att fortsätta. Telefonen stöds ej Avbryt  